module cpu(PC,INSTRUCTION,CLK,RESET);

endmodule